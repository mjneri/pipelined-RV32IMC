`timescale 1ns / 1ps

module if_id(

);

endmodule