`timescale 1ns / 1ps

module exe_mem(

);

endmodule