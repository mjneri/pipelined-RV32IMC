`timescale 1ns / 1ps

module storeblock(

);

endmodule