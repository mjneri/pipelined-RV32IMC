`timescale 1ns / 1ps

module BHT(
	input CLK,
	input nrst,

	
);


endmodule