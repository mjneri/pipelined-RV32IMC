`timescale 1ns / 1ps

module id_exe(

);

endmodule
