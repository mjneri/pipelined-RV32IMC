`timescale 1ns / 1ps

module tb_pipereg_mem_wb();

endmodule