`timescale 1ns / 1ps

module tb_pipereg_if_id();

endmodule