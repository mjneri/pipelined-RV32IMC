`ifndef CONST_VH		// Guard prevents header file from being included more than once
`define CONST_VH

`define INT_SIG_WIDTH 4

`define MEM_DEPTH 2048
`define MEM_WIDTH 16
`define WORD_WIDTH 32

`define PC_ADDR_BITS 12

`endif	// CONST_VH