`timescale 1ns / 1ps
/*

    Compressed Instruction Decoder

    This module implements the decoder that translates the 
    
    The decoder is separate and will be in the ID stage instead.

*/

module compressed_decoder(
    input clk,
    input nrst,
    input [11:0] inst,
    output [31:0] out_inst
    );

    

endmodule